`ifndef REG_BUS_DEFINES__SV
`define REG_BUS_DEFINES__SV

// bus properties
`define REG_BUS_AW   8
`define REG_BUS_DW   8
`define FIFO_AW      8
`define FIFO_DW      8

`endif // REG_BUS_DEFINES__SV