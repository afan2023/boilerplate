`ifndef REG_BUS_DEFINES__SV
`define REG_BUS_DEFINES__SV

// bus properties
`define REG_BUS_AW   5
`define REG_BUS_DW   16

`endif // REG_BUS_DEFINES__SV