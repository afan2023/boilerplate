`ifndef REG_BUS_SEQUENCER__SV
`define REG_BUS_SEQUENCER__SV

typedef uvm_sequencer #(reg_bus_transaction) reg_bus_sequencer;

`endif // REG_BUS_SEQUENCER__SV