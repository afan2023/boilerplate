`ifndef FIFO_RST_IF__SV
`define FIFO_RST_IF__SV

interface fifo_rst_if (input clk, input wclk, input rclk);

   logic rst_n ;
   
endinterface

`endif // FIFO_RST_IF__SV